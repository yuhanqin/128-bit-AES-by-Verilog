`timescale 10ns/1nsmodule aes();  //clk,reset_in,b0_in,b1_inreg rst_;reg [8:1] din;reg [2:1] cmd;reg clk=0;always clk=#1~clk;wire [8:1] dout;top i_uut(  .clk(clk),  .rst_(rst_),  .din(din),  .cmd(cmd),  .dout(dout),  .ok(ok),  .ready(ready));initial begin    $dumpfile("top.vcd");      $dumpvars(0, i_uut);   endinitial begin  din=8'b0;  cmd = 2'b0;  rst_ = 0;  #10;  rst_ = 1;  #10;  cmd = 2'b01;  din=8'h00;  #2;  din=8'h04;  #2;  din=8'h12;  #2;  din=8'h14;  #2;  din=8'h12;  #2;  din=8'h04;  #2;  din=8'h12;  #2;  din=8'h00;  #2;  din=8'h0c;  #2;  din=8'h00;  #2;  din=8'h13;  #2;  din=8'h11;  #2;  din=8'h08;  #2;  din=8'h23;  #2;  din=8'h19;  #2;  din=8'h19;  #10;  cmd = 2'b10;  din=8'h24;  #2;  din=8'h75;  #2;  din=8'ha2;  #2;  din=8'hb3;  #2;  din=8'h34;  #2;  din=8'h75;  #2;  din=8'h56;  #2;  din=8'h88;  #2;  din=8'h31;  #2;  din=8'he2;  #2;  din=8'h12;  #2;  din=8'h00;  #2;  din=8'h13;  #2;  din=8'haa;  #2;  din=8'h54;  #2;  din=8'h87;  #10;  cmd = 2'b11;  #100;    $finish();endendmodule